library ieee;
use ieee.std_logic_1164.all;

package memory_cell_pkg is

   constant memory_cell_parallelism_bit   : natural := 1;
   constant memory_cell_parallelism_delay : time    := 0 ns;

end package;
