----------------------------------------------------------------------------------
--! @file counter_modulo_n_pkg.vhd
--! @author Antonio Riccio
--! @brief Configuration values for the counter_modulo_n
--! @version 1.0
--! @date 30/07/2020
--! @copyright GNU Public License
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

package counter_modulo_n_pkg is

   constant counter_modulo : natural := 16;

end package;
