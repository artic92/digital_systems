library ieee;
use ieee.std_logic_1164.all;

package counter_modulo_n_pkg is

   constant counter_modulo : natural := 16;

end package;
