library ieee;
use ieee.std_logic_1164.all;

package register_n_bit_pkg is

   constant register_parallelism_bit   : natural := 1;
   constant register_parallelism_delay : time    := 0 ns;

end package;
